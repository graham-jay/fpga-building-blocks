module mux4 (

);

endmodule
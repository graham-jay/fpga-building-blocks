module dff (

);

endmodule
`include "../rtl/mux2.sv"

module mux2_tb ();
    

    mux2 DUT (

    );

    initial begin

    end

    task check_output(input reg value);

    endtask

endmodule

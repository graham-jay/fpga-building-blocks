`include "../rtl/dff.sv"

module dff_tb ();

    dff DUT (

    );

    initial begin

    end

    task check_output(input reg value);

    endtask

endmodule

`include "../rtl/mux4.sv"

module mux4_tb ();


    mux4 DUT (

    );

    initial begin

    end

    task check_output(input reg value);

    endtask

endmodule

module mux2 (

);

endmodule